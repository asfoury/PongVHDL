architecture rtl of movement_full is



begin


end architecture rtl;
