architecture rtl of pong is
begin

end architecture rtl; 
